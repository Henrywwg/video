module VGA();
    


endmodule
